module top (
    input               ext_clk_in,
    input               ext_rst_in,
    output     [03:00]  fpga_led
);


    assign fpga_led = 4'h0;

    zynq zynq (
        .DDR_addr                   (DDR_addr),
        .DDR_ba                     (DDR_ba),
        .DDR_cas_n                  (DDR_cas_n),
        .DDR_ck_n                   (DDR_ck_n),
        .DDR_ck_p                   (DDR_ck_p),
        .DDR_cke                    (DDR_cke),
        .DDR_cs_n                   (DDR_cs_n),
        .DDR_dm                     (DDR_dm),
        .DDR_dq                     (DDR_dq),
        .DDR_dqs_n                  (DDR_dqs_n),
        .DDR_dqs_p                  (DDR_dqs_p),
        .DDR_odt                    (DDR_odt),
        .DDR_ras_n                  (DDR_ras_n),
        .DDR_reset_n                (DDR_reset_n),
        .DDR_we_n                   (DDR_we_n),
        .ENET1_EXT_INTIN            (ENET1_EXT_INTIN),
        .FIXED_IO_ddr_vrn           (FIXED_IO_ddr_vrn),
        .FIXED_IO_ddr_vrp           (FIXED_IO_ddr_vrp),
        .FIXED_IO_mio               (FIXED_IO_mio),
        .FIXED_IO_ps_clk            (FIXED_IO_ps_clk),
        .FIXED_IO_ps_porb           (FIXED_IO_ps_porb),
        .FIXED_IO_ps_srstb          (FIXED_IO_ps_srstb),
        .GMII_ETHERNET_1_col        (GMII_ETHERNET_1_col),
        .GMII_ETHERNET_1_crs        (GMII_ETHERNET_1_crs),
        .GMII_ETHERNET_1_rx_clk     (GMII_ETHERNET_1_rx_clk),
        .GMII_ETHERNET_1_rx_dv      (GMII_ETHERNET_1_rx_dv),
        .GMII_ETHERNET_1_rx_er      (GMII_ETHERNET_1_rx_er),
        .GMII_ETHERNET_1_rxd        (GMII_ETHERNET_1_rxd),
        .GMII_ETHERNET_1_tx_clk     (GMII_ETHERNET_1_tx_clk),
        .GMII_ETHERNET_1_tx_en      (GMII_ETHERNET_1_tx_en),
        .GMII_ETHERNET_1_tx_er      (GMII_ETHERNET_1_tx_er),
        .GMII_ETHERNET_1_txd        (GMII_ETHERNET_1_txd),
        .IIC_0_scl_i                (IIC_0_scl_i),
        .IIC_0_scl_o                (IIC_0_scl_o),
        .IIC_0_scl_t                (IIC_0_scl_t),
        .IIC_0_sda_i                (IIC_0_sda_i),
        .IIC_0_sda_o                (IIC_0_sda_o),
        .IIC_0_sda_t                (IIC_0_sda_t),
        .M01_AXI_araddr             (M01_AXI_araddr),
        .M01_AXI_arprot             (M01_AXI_arprot),
        .M01_AXI_arready            (M01_AXI_arready),
        .M01_AXI_arvalid            (M01_AXI_arvalid),
        .M01_AXI_awaddr             (M01_AXI_awaddr),
        .M01_AXI_awprot             (M01_AXI_awprot),
        .M01_AXI_awready            (M01_AXI_awready),
        .M01_AXI_awvalid            (M01_AXI_awvalid),
        .M01_AXI_bready             (M01_AXI_bready),
        .M01_AXI_bresp              (M01_AXI_bresp),
        .M01_AXI_bvalid             (M01_AXI_bvalid),
        .M01_AXI_rdata              (M01_AXI_rdata),
        .M01_AXI_rready             (M01_AXI_rready),
        .M01_AXI_rresp              (M01_AXI_rresp),
        .M01_AXI_rvalid             (M01_AXI_rvalid),
        .M01_AXI_wdata              (M01_AXI_wdata),
        .M01_AXI_wready             (M01_AXI_wready),
        .M01_AXI_wstrb              (M01_AXI_wstrb),
        .M01_AXI_wvalid             (M01_AXI_wvalid),
        .M02_AXI_araddr             (M02_AXI_araddr),
        .M02_AXI_arprot             (M02_AXI_arprot),
        .M02_AXI_arready            (M02_AXI_arready),
        .M02_AXI_arvalid            (M02_AXI_arvalid),
        .M02_AXI_awaddr             (M02_AXI_awaddr),
        .M02_AXI_awprot             (M02_AXI_awprot),
        .M02_AXI_awready            (M02_AXI_awready),
        .M02_AXI_awvalid            (M02_AXI_awvalid),
        .M02_AXI_bready             (M02_AXI_bready),
        .M02_AXI_bresp              (M02_AXI_bresp),
        .M02_AXI_bvalid             (M02_AXI_bvalid),
        .M02_AXI_rdata              (M02_AXI_rdata),
        .M02_AXI_rready             (M02_AXI_rready),
        .M02_AXI_rresp              (M02_AXI_rresp),
        .M02_AXI_rvalid             (M02_AXI_rvalid),
        .M02_AXI_wdata              (M02_AXI_wdata),
        .M02_AXI_wready             (M02_AXI_wready),
        .M02_AXI_wstrb              (M02_AXI_wstrb),
        .M02_AXI_wvalid             (M02_AXI_wvalid),
        .M03_AXI_araddr             (M03_AXI_araddr),
        .M03_AXI_arprot             (M03_AXI_arprot),
        .M03_AXI_arready            (M03_AXI_arready),
        .M03_AXI_arvalid            (M03_AXI_arvalid),
        .M03_AXI_awaddr             (M03_AXI_awaddr),
        .M03_AXI_awprot             (M03_AXI_awprot),
        .M03_AXI_awready            (M03_AXI_awready),
        .M03_AXI_awvalid            (M03_AXI_awvalid),
        .M03_AXI_bready             (M03_AXI_bready),
        .M03_AXI_bresp              (M03_AXI_bresp),
        .M03_AXI_bvalid             (M03_AXI_bvalid),
        .M03_AXI_rdata              (M03_AXI_rdata),
        .M03_AXI_rready             (M03_AXI_rready),
        .M03_AXI_rresp              (M03_AXI_rresp),
        .M03_AXI_rvalid             (M03_AXI_rvalid),
        .M03_AXI_wdata              (M03_AXI_wdata),
        .M03_AXI_wready             (M03_AXI_wready),
        .M03_AXI_wstrb              (M03_AXI_wstrb),
        .M03_AXI_wvalid             (M03_AXI_wvalid),
        .MDIO_ETHERNET_1_mdc        (MDIO_ETHERNET_1_mdc),
        .MDIO_ETHERNET_1_mdio_i     (MDIO_ETHERNET_1_mdio_i),
        .MDIO_ETHERNET_1_mdio_o     (MDIO_ETHERNET_1_mdio_o),
        .MDIO_ETHERNET_1_mdio_t     (MDIO_ETHERNET_1_mdio_t),
        .USBIND_0_port_indctl       (USBIND_0_port_indctl),
        .USBIND_0_vbus_pwrfault     (USBIND_0_vbus_pwrfault),
        .USBIND_0_vbus_pwrselect    (USBIND_0_vbus_pwrselect),
        .cpu_if_araddr              (cpu_if_araddr),
        .cpu_if_arprot              (cpu_if_arprot),
        .cpu_if_arready             (cpu_if_arready),
        .cpu_if_arvalid             (cpu_if_arvalid),
        .cpu_if_awaddr              (cpu_if_awaddr),
        .cpu_if_awprot              (cpu_if_awprot),
        .cpu_if_awready             (cpu_if_awready),
        .cpu_if_awvalid             (cpu_if_awvalid),
        .cpu_if_bready              (cpu_if_bready),
        .cpu_if_bresp               (cpu_if_bresp),
        .cpu_if_bvalid              (cpu_if_bvalid),
        .cpu_if_rdata               (cpu_if_rdata),
        .cpu_if_rready              (cpu_if_rready),
        .cpu_if_rresp               (cpu_if_rresp),
        .cpu_if_rvalid              (cpu_if_rvalid),
        .cpu_if_wdata               (cpu_if_wdata),
        .cpu_if_wready              (cpu_if_wready),
        .cpu_if_wstrb               (cpu_if_wstrb),
        .cpu_if_wvalid              (cpu_if_wvalid),
        .zynq_clk                   (zynq_clk),
        .zynq_resetn                (zynq_resetn)
    );

    mb_sys mb_sys (
        .mb_clk_in          ( mb_clk_in     ),
        .mb_rst_n_in        ( 1'b1          ) 
    );

    

endmodule